module AGDC_moore_tb ();

 reg UP_Max_tb , Activate_tb , DN_Max_tb ;
 reg CLK_tb , RST_tb ;
 wire UP_M_tb , DN_M_tb ;

parameter clk_p = 20 ;

always 
 begin
  #(clk_p/2) CLK_tb = ~CLK_tb ;
 end

AGDC_moore dut (.UP_Max(UP_Max_tb) , 
            .Activate(Activate_tb) , 
            .DN_Max(DN_Max_tb) , 
            .CLK(CLK_tb) , 
            .RST(RST_tb) , 
            .UP_M(UP_M_tb) , 
            .DN_M(DN_M_tb)) ;

task initialize ;
 begin
  UP_Max_tb = 1'b0 ;
  Activate_tb = 1'b0 ;
  DN_Max_tb = 1'b0 ;
  CLK_tb = 1'b0 ;
 end
 endtask 

task reset ;
 begin
  RST_tb = 1'b1 ;
  #clk_p 
  RST_tb = 1'b0 ;
  #clk_p 
  RST_tb = 1'b1 ;
 end
 endtask
initial 
 begin
  initialize () ;
  reset () ;
 
 
if ((UP_M_tb == 1'b0) && (DN_M_tb == 1'b0))
 $display (" reset case passed ") ;
else
 $display (" reset case failed ") ;

Activate_tb = 1'b1 ;
UP_Max_tb = 1'b1 ;

#clk_p 

if ((UP_M_tb == 1'b0) && (DN_M_tb == 1'b1))
 $display (" UP case passed ") ;
else
 $display (" UP case failed ") ;

DN_Max_tb = 1'b1 ;

#clk_p

if ((UP_M_tb == 1'b0) && (DN_M_tb == 1'b0))
 $display (" ideal case passed ") ;
else
 $display (" ideal case failed ") ;

UP_Max_tb = 1'b0 ;

#clk_p

if ((UP_M_tb == 1'b1) && (DN_M_tb == 1'b0))
 $display (" DN case passed ") ;
else
 $display (" DN case failed ") ;

end

endmodule