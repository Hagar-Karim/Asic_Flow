module ALU_16B 
(
  input wire [15:0] A , B ,
  input wire [3:0]  ALU_FUN ,
  input wire clk ,
  output reg [15:0] ALU_OUT ,
  output reg Carry_Flag ,
  output reg Arith_Flag ,
  output reg Logic_Flag ,
  output reg CMP_Flag ,
  output reg Shift_Flag

);

always@ (posedge clk)
 begin
   case(ALU_FUN)
    
    4'b0000 : 
    begin 
    {Carry_Flag , ALU_OUT} <= A + B ;
     Arith_Flag <= 1'b1;
     Logic_Flag <= 1'b0;
     CMP_Flag <= 1'b0 ;
     Shift_Flag <= 1'b0 ;
    end
    4'b0001 :
    begin
    {Carry_Flag , ALU_OUT} <= A - B ;
     Arith_Flag <= 1'b1;
     Logic_Flag <= 1'b0;
     CMP_Flag <= 1'b0 ;
     Shift_Flag <= 1'b0 ;
    end
    4'b0010 :
    begin
    ALU_OUT <= A * B ;
    Arith_Flag <= 1'b1;
    Logic_Flag <= 1'b0;
    CMP_Flag <= 1'b0 ;
    Shift_Flag <= 1'b0 ;
    Carry_Flag <= 1'b0 ;
    end
    4'b0011 :
    begin
    ALU_OUT <= A / B ;
    Arith_Flag <= 1'b1;
    Logic_Flag <= 1'b0;
    CMP_Flag <= 1'b0 ;
    Shift_Flag <= 1'b0 ;
    Carry_Flag <= 1'b0 ;
    end
    4'b0100 :
    begin
    ALU_OUT <= A & B ;
    Arith_Flag <= 1'b0 ;
    Logic_Flag <= 1'b1 ;
    CMP_Flag <= 1'b0 ;
    Shift_Flag <= 1'b0 ;
    Carry_Flag <= 1'b0 ;
    end
    4'b0101 :
     begin
      ALU_OUT <= A | B ;
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b1 ;
      CMP_Flag <= 1'b0 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b0110 :
     begin
      ALU_OUT <= ~(A & B) ;
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b1 ;
      CMP_Flag <= 1'b0 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b0111 :
     begin
      ALU_OUT <= ~(A | B) ;
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b1 ;
      CMP_Flag <= 1'b0 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b1000 :
     begin
      ALU_OUT <= A ^ B ;
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b1 ;
      CMP_Flag <= 1'b0 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b1001 :
     begin
      ALU_OUT <= ~(A ^ B) ;
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b1 ;
      CMP_Flag <= 1'b0 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b1010 :
     begin
      if (A == B)
       ALU_OUT <= 16'b1 ;
      else
       ALU_OUT <= 1'b0 ;

      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b0 ;
      CMP_Flag <= 1'b1 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b1011 :
     begin
      if (A > B)
       ALU_OUT <= 16'b10 ;
      else
       ALU_OUT <= 1'b0 ;
       
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b0 ;
      CMP_Flag <= 1'b1 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b1100 :
     begin
      if (A < B)
       ALU_OUT <= 16'b11 ;
      else
       ALU_OUT <= 1'b0 ;
       
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b0 ;
      CMP_Flag <= 1'b1 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b1101 :
     begin
      ALU_OUT <= A >> 1 ;
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b0 ;
      CMP_Flag <= 1'b0 ;
      Shift_Flag <= 1'b1 ;
      Carry_Flag <= 1'b0 ;
    end
    4'b1110 :
     begin
      ALU_OUT <= A << 1 ;
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b0 ;
      CMP_Flag <= 1'b0 ;
      Shift_Flag <= 1'b1 ;
      Carry_Flag <= 1'b0 ;
    end
   default :
   begin
      ALU_OUT <= 1'b0 ;
      Arith_Flag <= 1'b0 ;
      Logic_Flag <= 1'b0 ;
      CMP_Flag <= 1'b0 ;
      Shift_Flag <= 1'b0 ;
      Carry_Flag <= 1'b0 ;
    end

  endcase
 end
 endmodule